-- FILEPATH: /pipe/DF_EX.vhd

library ieee;
use ieee.std_logic_1164.all;

entity DF_MEM is
  port (
    -- Adicione aqui as portas de entrada e saída do componente
  );
end entity DF_MEM;

architecture rtl of DF_MEM is
begin
  -- Adicione aqui a lógica do componente
end architecture rtl;
