------------------------------------------------------
--! @file ALU.vhdl
--! @brief Testbench for my very own ALU!
--! @author Miguel Aguena (miguel.aguena@usp.br)
--! @date 2021-11-08
-------------------------------------------------------

entity tb is
end tb;
    
    architecture testbench_1 of tb is
        component rom is
            port (
                addr : in  bit_vector(7 downto 0);
                data : out bit_vector(31 downto 0)
            );
        end component rom;
        component polilegsc is
            port (
                clock, reset : in bit;
                --Data Memory
                dmem_addr : out bit_vector(63 downto 0);
                dmem_dati : out bit_vector(63 downto 0);
                dmem_dato : in bit_vector(63 downto 0);
                dmem_we : out bit;
                --Instruction Memory
                imem_addr : out bit_vector(63 downto 0);
                imem_data : in bit_vector(31 downto 0)
            );
        end component polilegsc;
        component ram is
            generic (
                addr_s : natural := 8;
                word_s : natural := 64;
                a : natural := 32;
                b : natural := 96
            );
            port (
                ck     : in  bit;
                rd, wr : in  bit;
                addr   : in  bit_vector(addr_s-1 downto 0);
                data_i : in  bit_vector(word_s-1 downto 0);
                data_o : out bit_vector(word_s-1 downto 0)
            );
        end component ram;
    
        signal imem_addr_aux : bit_vector(63 downto 0);
        signal imem_data_aux : bit_vector(31 downto 0);
        signal dmem_addr_aux : bit_vector(63 downto 0);
        signal dmem_dati_aux : bit_vector(63 downto 0);
        signal dmem_dato_aux : bit_vector(63 downto 0);
        signal dmem_we_aux : bit;
        signal clock : bit;
    begin
        ROM_INSTR: rom port map (
            addr => imem_addr_aux(7 downto 0),
            data => imem_data_aux
        );

        POLILEG_CPU: polilegsc port map (
            clock => clock,
            reset => '0',
            --Data Memory
            dmem_addr => dmem_addr_aux,
            dmem_dati => dmem_dati_aux,
            dmem_dato => dmem_dato_aux,
            dmem_we => dmem_we_aux,
            --Instruction Memory
            imem_addr => imem_addr_aux,
            imem_data => imem_data_aux
        );

        RAM_DATA: ram generic map (8, 64, 63, 56) port map (
            ck => clock,
            rd => '1',
            wr => dmem_we_aux,
            addr => dmem_addr_aux(7 downto 0),
            data_i => dmem_dati_aux,
            data_o => dmem_dato_aux
        );
    
        p: process is
            type pattern_type is record
                clock : bit;
                a : bit;
            end record;
    
            type pattern_array is array (natural range <>) of pattern_type;
            constant patterns : pattern_array := (
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0'),
                ('1', '0'),
                ('0', '0')
            );
        begin
            for k in patterns'range loop
                clock <= patterns(k).clock;
    
                wait for 1 ns;
            end loop;
    
            assert false report "end of test" severity note;
            wait;
        end process;
    end architecture testbench_1;